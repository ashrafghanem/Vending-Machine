----------------------------------------------------------------------------------
-- COMPANY: 
-- ENGINEER: 
-- 
-- CREATE DATE:    19:34:17 11/30/2017 
-- DESIGN NAME: 
-- MODULE NAME:    VENDINGMACHINE - BEHAVIORAL 
-- PROJECT NAME: 
-- TARGET DEVICES: 
-- TOOL VERSIONS: 
-- DESCRIPTION: 
--
-- DEPENDENCIES: 
--
-- REVISION: 
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF INSTANTIATING
-- ANY XILINX PRIMITIVES IN THIS CODE.
--LIBRARY UNISIM;
--USE UNISIM.VCOMPONENTS.ALL;

ENTITY VENDINGMACHINE IS
	PORT( S,CLOCK,RESET: IN STD_LOGIC;
			C: IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
			P: IN  STD_LOGIC_VECTOR(2 DOWNTO 1);
			R: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			PRODUCT: OUT STD_LOGIC_VECTOR(2 DOWNTO 1));
END VENDINGMACHINE;

ARCHITECTURE BEHAVIORAL OF VENDINGMACHINE IS
		TYPE STATE IS (S0,S1,S2,S3);
		SIGNAL CURR_STATE: STATE := S0;
		SIGNAL NEXT_STATE: STATE ;
		
		SIGNAL SUM,PRICE: INTEGER RANGE 0 TO 9:= 0;		
		
BEGIN
		CLOCKED: PROCESS (RESET, CLOCK)
		BEGIN
			IF(RESET='1') THEN
				CURR_STATE <= S0;
			ELSIF (CLOCK 'EVENT AND CLOCK='1') THEN
				IF CURR_STATE = S1 THEN
					SUM <= 0;
					PRICE <= 0;
					PRODUCT <= "00";
					R <= "000";
					IF (P(1) = '1') THEN
						PRICE <= 6;
					ELSIF (P(2) = '1') THEN
						PRICE <= 5;
					END IF;
					
				ELSIF CURR_STATE = S2 THEN
					IF(SUM < PRICE) THEN
						IF    (C(0) = '1') THEN SUM <= SUM + 1;
						ELSIF (C(1) = '1') THEN SUM <= SUM + 2;
						ELSIF (C(2) = '1') THEN SUM <= SUM + 4;
						END IF;
					ELSE
						IF (P(2)='1') THEN PRODUCT(2)<='1';
						ELSE PRODUCT(1)<='1';
						END IF;
					END IF;
					
				ELSIF CURR_STATE = S3 THEN
					IF    (SUM-PRICE=3) THEN R <= "011";
					ELSIF (SUM-PRICE=2) THEN R <= "010";
					ELSIF (SUM-PRICE=1) THEN R <= "001";
					END IF;
				END IF;
			CURR_STATE <= NEXT_STATE;
			END IF;
		END PROCESS CLOCKED;
		
		COMBINATIONAL: PROCESS(CURR_STATE,S,C,P)
		BEGIN
			CASE CURR_STATE IS
				WHEN S0 => 
					IF S='1' THEN 
						NEXT_STATE <= S1;
					ELSE
						NEXT_STATE <= S0;
					END IF;
				WHEN S1 =>
					IF P(1)='1' THEN
						NEXT_STATE <= S2;
					ELSE
						IF P(2) = '1' THEN
							NEXT_STATE <= S2;
						ELSE
							NEXT_STATE <= S1;
						END IF;
					END IF;
				WHEN S2 =>
					IF SUM < PRICE THEN
						NEXT_STATE <= S2;
					ELSE
						NEXT_STATE <= S3;
					END IF;
				WHEN S3 =>
					NEXT_STATE <= S0;
				WHEN OTHERS =>
					NEXT_STATE <= S0;
			END CASE;
		END PROCESS COMBINATIONAL;
			
END BEHAVIORAL;

